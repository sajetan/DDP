`timescale 1ns / 1ps

module montgomery(
    input          clk,
    input          resetn,
    input          start,
    input  [511:0] in_a,
    input  [511:0] in_b,
    input  [511:0] in_m,
    output [511:0] result,  
    output         done
     );
 
    
    // Student tasks:
    // 1. Instantiate an Adder
    // 2. Use the Adder to implement the Montgomery multiplier in hardware.
    // 3. Use tb_montgomery.v to simulate your design.
    
    
    // This always block was added to ensure the tool doesn't trim away the montgomery module.
    // Feel free to remove this block
    reg [511:0] r_result;
    always @(posedge(clk))
    begin
        r_result <= {512{1'b1}};
    end
    assign result = r_result;

    assign done = 1;
endmodule